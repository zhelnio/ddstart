
module top
(
    input  io_72,
    input  io_73,
    output io_74
);
    assign io_74 = io_72 ^ io_73;

endmodule
